library IEEE ;
use IEEE.STD_LOGIC_1164.all ;

package	constants is
	type TPicoType is ( pbtI, pbtII, pbt3, pbtS ) ;
	constant PicoType : TPicoType := pbt3 ;
	function ADDRSIZE return natural ;
	function INSTSIZE return natural ;
	function JADDRSIZE return natural ;
	function JDATASIZE return natural ;
end package ;

package body constants is
	function ADDRSIZE return natural is
	begin
		case PicoType is
		when pbtI => return 8 ;
		when pbtII => return 10 ;
		when pbt3 => return 10 ;
		when pbtS => return 10 ;
		end case ;
	end ;
	function INSTSIZE return natural is 
	begin
		case PicoType is
		when pbtI => return 16 ;
		when pbtII => return 18 ;
		when pbt3 => return 18 ;
		when pbtS => return 18 ;
		end case ;
	end ;
	function JADDRSIZE return natural is
	begin
		case PicoType is
		when pbtI => return 9 ;
		when pbtII => return 11 ;
		when pbt3 => return 11 ;
		when pbtS => return 10 ;
		end case ;
	end ;
	function JDATASIZE return natural is
	begin
		case PicoType is
		when pbtI => return 8 ;
		when pbtII => return 9 ;
		when pbt3 => return 9 ;
		when pbtS => return 20 ;
		end case ;
	end ;
end package body ;


library IEEE ;
use IEEE.STD_LOGIC_1164.all ;
use IEEE.STD_LOGIC_ARITH.all ;
use IEEE.STD_LOGIC_UNSIGNED.all ;

library unisim ;
use unisim.vcomponents.all ;

use constants.all;

entity prog_rom is
    port ( 
        clk : in std_logic ;
        reset : out std_logic ;
        address : in std_logic_vector( ADDRSIZE - 1 downto 0 ) ;
        instruction : out std_logic_vector( INSTSIZE - 1 downto 0 )
    ) ;
end entity prog_rom ;

architecture mix of prog_rom is
    component jtag_shifter is
        port ( 
			clk : in std_logic ;
			user1 : out std_logic ;
            write : out std_logic ;
            addr : out std_logic_vector( JADDRSIZE - 1 downto 0 ) ;
            data : out std_logic_vector( JDATASIZE - 1 downto 0 )
        ) ;
    end component ;

    signal jaddr : std_logic_vector( JADDRSIZE - 1 downto 0 ) ;
    signal jdata : std_logic_vector( JDATASIZE - 1 downto 0 ) ;
    signal juser1 : std_logic ;
    signal jwrite : std_logic ;

    attribute INIT_00 : string ;
    attribute INIT_01 : string ;
    attribute INIT_02 : string ;
    attribute INIT_03 : string ;
    attribute INIT_04 : string ;
    attribute INIT_05 : string ;
    attribute INIT_06 : string ;
    attribute INIT_07 : string ;
    attribute INIT_08 : string ;
    attribute INIT_09 : string ;
    attribute INIT_0A : string ;
    attribute INIT_0B : string ;
    attribute INIT_0C : string ;
    attribute INIT_0D : string ;
    attribute INIT_0E : string ;
    attribute INIT_0F : string ;
    attribute INIT_10 : string ;
    attribute INIT_11 : string ;
    attribute INIT_12 : string ;
    attribute INIT_13 : string ;
    attribute INIT_14 : string ;
    attribute INIT_15 : string ;
    attribute INIT_16 : string ;
    attribute INIT_17 : string ;
    attribute INIT_18 : string ;
    attribute INIT_19 : string ;
    attribute INIT_1A : string ;
    attribute INIT_1B : string ;
    attribute INIT_1C : string ;
    attribute INIT_1D : string ;
    attribute INIT_1E : string ;
    attribute INIT_1F : string ;
    attribute INIT_20 : string ;
    attribute INIT_21 : string ;
    attribute INIT_22 : string ;
    attribute INIT_23 : string ;
    attribute INIT_24 : string ;
    attribute INIT_25 : string ;
    attribute INIT_26 : string ;
    attribute INIT_27 : string ;
    attribute INIT_28 : string ;
    attribute INIT_29 : string ;
    attribute INIT_2A : string ;
    attribute INIT_2B : string ;
    attribute INIT_2C : string ;
    attribute INIT_2D : string ;
    attribute INIT_2E : string ;
    attribute INIT_2F : string ;
    attribute INIT_30 : string ;
    attribute INIT_31 : string ;
    attribute INIT_32 : string ;
    attribute INIT_33 : string ;
    attribute INIT_34 : string ;
    attribute INIT_35 : string ;
    attribute INIT_36 : string ;
    attribute INIT_37 : string ;
    attribute INIT_38 : string ;
    attribute INIT_39 : string ;
    attribute INIT_3A : string ;
    attribute INIT_3B : string ;
    attribute INIT_3C : string ;
    attribute INIT_3D : string ;
    attribute INIT_3E : string ;
    attribute INIT_3F : string ;
    attribute INITP_00 : string ;
    attribute INITP_01 : string ;
    attribute INITP_02 : string ;
    attribute INITP_03 : string ;
    attribute INITP_04 : string ;
    attribute INITP_05 : string ;
    attribute INITP_06 : string ;
    attribute INITP_07 : string ;
begin
	I18 : if (PicoType = pbtII) or (PicoType = pbt3) generate
	    attribute INIT_00 of bram : label is "40FE502B40FFB0002F40A0000D00CF40AF04540B40FD40F01000C0F04001C001" ;
	    attribute INIT_01 of bram : label is "CF01A000AF04501F400050204001542D2DFF54232F20AF7F80FD50152F80502F" ;
	    attribute INIT_02 of bram : label is "2CFFA000AF04A000CF80404F03E0A0008D01F0D05C294D20FC00A0001C00CF20" ;
	    attribute INIT_03 of bram : label is "50DE400E50AA400450974003507C400250704001505F4000600003E0544F03E1" ;
	    attribute INIT_04 of bram : label is "2F0103E2514D400C505E400D5141400B512D400A50EE40095124400850E5400F" ;
	    attribute INIT_05 of bram : label is "4D044000A000AF04C3F15458240144F203FEC3F15453240144F2E3FFC3F1B400" ;
	    attribute INIT_06 of bram : label is "404F03DA5468CD0182018001D3207300584F941003E314206201CD030002584F" ;
	    attribute INIT_07 of bram : label is "62010002584F4D05404F03DA5475CD018001D32073006201CD030002584F4D04" ;
	    attribute INIT_08 of bram : label is "7300C2018001D32073008201584F941003E31420544F2D01CD03544F220103E5" ;
	    attribute INIT_09 of bram : label is "504F20FF03E360026101544F4D04B4002F01404F03DA548BCD0282038001D320" ;
	    attribute INIT_0A of bram : label is "60026101544F4D04B4002F0140B554A4C001810100C0531000D7584F92101200" ;
	    attribute INIT_0B of bram : label is "A000AF04C3F154BA240144F203FE00C013C0B4002F0154B1C00100C0531000D7" ;
	    attribute INIT_0C of bram : label is "CE01041E5CD38E01C3F154C8240144F203FFC5FD153058C843FDFC30B4002F01" ;
	    attribute INIT_0D of bram : label is "000400D7A000C3F103FD0E000C00B4002F0140C81350B40043FF54CFC40154CF" ;
	    attribute INIT_0E of bram : label is "1980680140B554E8CD01800100C07300CD01000000D740B554E0C00100C00308" ;
	    attribute INIT_0F of bram : label is "03E7550149C05117A9C054F7C60107000806544F03E658F7481007000604A83F" ;
	    attribute INIT_10 of bram : label is "012AB12090300121550F4980610360021B701A80544F03E051064D02CD03544F" ;
	    attribute INIT_11 of bram : label is "00C0132000C0012100D7544F03E0511B4D03115010405D17012A115010405913" ;
	    attribute INIT_12 of bram : label is "2F04584F4D05A000F310D200404F03DADF00AFFBA0046001A000A700880440B5" ;
	    attribute INIT_13 of bram : label is "03DA553CCD018001544F24F803E3A40093D01320141062026101CD04000350FF" ;
	    attribute INIT_14 of bram : label is "4D04B4002F0140B55549C00100C000D7600362026101544F4D05B4002F01404F" ;
	    attribute INIT_15 of bram : label is "00000000000000008001000240B55554C001810100C0731000D760026101544F" ;
	    attribute INIT_16 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_17 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_18 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_19 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1A of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1F of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_20 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_21 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_22 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_23 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_24 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_25 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_26 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_27 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_28 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_29 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2A of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2F of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_30 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_31 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_32 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_33 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_34 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_35 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_36 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_37 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_38 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_39 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3A of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3F of bram : label is "415A000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_00 of bram : label is "0DCD604DCD58D01378B42D0A4DDDDDDDDDDDDD0C62326D20237774777660342F" ;
	    attribute INITP_01 of bram : label is "3736B3400F5C4FDC3A0272774DB413498B4327730D9F5CF4D0367356161D0D74" ;
	    attribute INITP_02 of bram : label is "000000000000000000FF5CC367DF036735D14013765C0097CFF343C3D7D00CD7" ;
	    attribute INITP_03 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_04 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_05 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_06 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_07 of bram : label is "C000000000000000000000000000000000000000000000000000000000000000" ;
	begin
	    bram : component RAMB16_S9_S18
	        generic map (
	            INIT_00 => X"40FE502B40FFB0002F40A0000D00CF40AF04540B40FD40F01000C0F04001C001",
	            INIT_01 => X"CF01A000AF04501F400050204001542D2DFF54232F20AF7F80FD50152F80502F",
	            INIT_02 => X"2CFFA000AF04A000CF80404F03E0A0008D01F0D05C294D20FC00A0001C00CF20",
	            INIT_03 => X"50DE400E50AA400450974003507C400250704001505F4000600003E0544F03E1",
	            INIT_04 => X"2F0103E2514D400C505E400D5141400B512D400A50EE40095124400850E5400F",
	            INIT_05 => X"4D044000A000AF04C3F15458240144F203FEC3F15453240144F2E3FFC3F1B400",
	            INIT_06 => X"404F03DA5468CD0182018001D3207300584F941003E314206201CD030002584F",
	            INIT_07 => X"62010002584F4D05404F03DA5475CD018001D32073006201CD030002584F4D04",
	            INIT_08 => X"7300C2018001D32073008201584F941003E31420544F2D01CD03544F220103E5",
	            INIT_09 => X"504F20FF03E360026101544F4D04B4002F01404F03DA548BCD0282038001D320",
	            INIT_0A => X"60026101544F4D04B4002F0140B554A4C001810100C0531000D7584F92101200",
	            INIT_0B => X"A000AF04C3F154BA240144F203FE00C013C0B4002F0154B1C00100C0531000D7",
	            INIT_0C => X"CE01041E5CD38E01C3F154C8240144F203FFC5FD153058C843FDFC30B4002F01",
	            INIT_0D => X"000400D7A000C3F103FD0E000C00B4002F0140C81350B40043FF54CFC40154CF",
	            INIT_0E => X"1980680140B554E8CD01800100C07300CD01000000D740B554E0C00100C00308",
	            INIT_0F => X"03E7550149C05117A9C054F7C60107000806544F03E658F7481007000604A83F",
	            INIT_10 => X"012AB12090300121550F4980610360021B701A80544F03E051064D02CD03544F",
	            INIT_11 => X"00C0132000C0012100D7544F03E0511B4D03115010405D17012A115010405913",
	            INIT_12 => X"2F04584F4D05A000F310D200404F03DADF00AFFBA0046001A000A700880440B5",
	            INIT_13 => X"03DA553CCD018001544F24F803E3A40093D01320141062026101CD04000350FF",
	            INIT_14 => X"4D04B4002F0140B55549C00100C000D7600362026101544F4D05B4002F01404F",
	            INIT_15 => X"00000000000000008001000240B55554C001810100C0731000D760026101544F",
	            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3F => X"415A000000000000000000000000000000000000000000000000000000000000",
	            INITP_00 => X"0DCD604DCD58D01378B42D0A4DDDDDDDDDDDDD0C62326D20237774777660342F",
	            INITP_01 => X"3736B3400F5C4FDC3A0272774DB413498B4327730D9F5CF4D0367356161D0D74",
	            INITP_02 => X"000000000000000000FF5CC367DF036735D14013765C0097CFF343C3D7D00CD7",
	            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_07 => X"C000000000000000000000000000000000000000000000000000000000000000"
	        )
	        port map (
	            DIB => "0000000000000000",
	            DIPB => "00",
	            ENB => '1',
	            WEB => '0',
	            SSRB => '0',
	            CLKB => clk,
	            ADDRB => address,
	            DOB => instruction( INSTSIZE - 3 downto 0 ),
	            DOPB => instruction( INSTSIZE - 1 downto INSTSIZE - 2 ),
	            DIA => jdata( JDATASIZE - 2 downto 0 ),
	            DIPA => jdata( JDATASIZE - 1 downto JDATASIZE - 1 ),
	            ENA => juser1,
	            WEA => jwrite,
	            SSRA => '0',
	            CLKA => clk,
	            ADDRA => jaddr,
	            DOA => open,
	            DOPA => open 
	        ) ;
	end generate ;

	I16 : if PicoType = pbtI generate
		attribute INIT_00 of bram : label is "40FE502B40FFB0002F40A0000D00CF40AF04540B40FD40F01000C0F04001C001" ;
		attribute INIT_01 of bram : label is "CF01A000AF04501F400050204001542D2DFF54232F20AF7F80FD50152F80502F" ;
		attribute INIT_02 of bram : label is "2CFFA000AF04A000CF80404F03E0A0008D01F0D05C294D20FC00A0001C00CF20" ;
		attribute INIT_03 of bram : label is "50DE400E50AA400450974003507C400250704001505F4000600003E0544F03E1" ;
		attribute INIT_04 of bram : label is "2F0103E2514D400C505E400D5141400B512D400A50EE40095124400850E5400F" ;
		attribute INIT_05 of bram : label is "4D044000A000AF04C3F15458240144F203FEC3F15453240144F2E3FFC3F1B400" ;
		attribute INIT_06 of bram : label is "404F03DA5468CD0182018001D3207300584F941003E314206201CD030002584F" ;
		attribute INIT_07 of bram : label is "62010002584F4D05404F03DA5475CD018001D32073006201CD030002584F4D04" ;
		attribute INIT_08 of bram : label is "7300C2018001D32073008201584F941003E31420544F2D01CD03544F220103E5" ;
		attribute INIT_09 of bram : label is "504F20FF03E360026101544F4D04B4002F01404F03DA548BCD0282038001D320" ;
		attribute INIT_0A of bram : label is "60026101544F4D04B4002F0140B554A4C001810100C0531000D7584F92101200" ;
		attribute INIT_0B of bram : label is "A000AF04C3F154BA240144F203FE00C013C0B4002F0154B1C00100C0531000D7" ;
		attribute INIT_0C of bram : label is "CE01041E5CD38E01C3F154C8240144F203FFC5FD153058C843FDFC30B4002F01" ;
		attribute INIT_0D of bram : label is "000400D7A000C3F103FD0E000C00B4002F0140C81350B40043FF54CFC40154CF" ;
		attribute INIT_0E of bram : label is "1980680140B554E8CD01800100C07300CD01000000D740B554E0C00100C00308" ;
		attribute INIT_0F of bram : label is "03E7550149C05117A9C054F7C60107000806544F03E658F7481007000604A83F" ;
	begin
	    bram : component RAMB4_S8_S16
	        generic map (
	            INIT_00 => X"40FE502B40FFB0002F40A0000D00CF40AF04540B40FD40F01000C0F04001C001",
	            INIT_01 => X"CF01A000AF04501F400050204001542D2DFF54232F20AF7F80FD50152F80502F",
	            INIT_02 => X"2CFFA000AF04A000CF80404F03E0A0008D01F0D05C294D20FC00A0001C00CF20",
	            INIT_03 => X"50DE400E50AA400450974003507C400250704001505F4000600003E0544F03E1",
	            INIT_04 => X"2F0103E2514D400C505E400D5141400B512D400A50EE40095124400850E5400F",
	            INIT_05 => X"4D044000A000AF04C3F15458240144F203FEC3F15453240144F2E3FFC3F1B400",
	            INIT_06 => X"404F03DA5468CD0182018001D3207300584F941003E314206201CD030002584F",
	            INIT_07 => X"62010002584F4D05404F03DA5475CD018001D32073006201CD030002584F4D04",
	            INIT_08 => X"7300C2018001D32073008201584F941003E31420544F2D01CD03544F220103E5",
	            INIT_09 => X"504F20FF03E360026101544F4D04B4002F01404F03DA548BCD0282038001D320",
	            INIT_0A => X"60026101544F4D04B4002F0140B554A4C001810100C0531000D7584F92101200",
	            INIT_0B => X"A000AF04C3F154BA240144F203FE00C013C0B4002F0154B1C00100C0531000D7",
	            INIT_0C => X"CE01041E5CD38E01C3F154C8240144F203FFC5FD153058C843FDFC30B4002F01",
	            INIT_0D => X"000400D7A000C3F103FD0E000C00B4002F0140C81350B40043FF54CFC40154CF",
	            INIT_0E => X"1980680140B554E8CD01800100C07300CD01000000D740B554E0C00100C00308",
	            INIT_0F => X"03E7550149C05117A9C054F7C60107000806544F03E658F7481007000604A83F"
	        )
			port map (
				DIB => "0000000000000000",  
				ENB => '1', 
				WEB => '0',
				RSTB =>	'0',
				CLKB => clk,
				ADDRB => address,
				DOB => instruction( INSTSIZE - 1 downto 0 ),  
				DIA => jdata( JDATASIZE - 1 downto 0 ),   
				ENA => juser1, 
				WEA => jwrite,
				RSTA => '0',
				CLKA => clk,
				ADDRA => jaddr,
				DOA => open  
			) ; 
	end generate ;

	I20 : if PicoType = pbtS generate
		attribute INIT_00 of ram_1 : label is "3131313131310030120203021231020002031313131013131312120003100233" ;
		attribute INIT_01 of ram_1 : label is "0031303112001031303111203100010313202310023100221031313131313131" ;
		attribute INIT_02 of ram_1 : label is "2023100302131303003121331130331031000312130311120112013100311310" ;
		attribute INIT_03 of ram_1 : label is "0313031223031000003311301033313003220002130213131031231001031021" ;
		attribute INIT_04 of ram_1 : label is "0311310110000103131211300000211330333303100330033113310000303113" ;
		attribute INIT_05 of ram_1 : label is "0000000000000000000000000000000000003333113030031213313300031213" ;
		attribute INIT_06 of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_07 of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_08 of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_09 of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0A of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0B of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0C of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0D of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0E of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0F of ram_1 : label is "3000000000000000000000000000000000000000000000000000000000000000" ;

		attribute INIT_00 of ram_2 : label is "54545454545460502AAAC40A8F54FA1CCAA54545252A8525454B2A0CA5441C4C" ;
		attribute INIT_01 of ram_2 : label is "6054405C8D76C054405C88D759016C0544AAC5240C524ECB2054545454545454" ;
		attribute INIT_02 of ram_2 : label is "AAC524001B25C0506654B245C80505915206654B2405C88D7C8D78590152C520" ;
		attribute INIT_03 of ram_2 : label is "0545A5C00505400A1645C807C0045C0000AC000B241B45C5C058C5240C154FB2" ;
		attribute INIT_04 of ram_2 : label is "05C8520A91166C05254AFD40DAA6AA8401000505411501150B905466115054C5" ;
		attribute INIT_05 of ram_2 : label is "0000000000000000000000000000000000008045C80706654B245C0066654B24" ;
		attribute INIT_06 of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_07 of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_08 of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_09 of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0A of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0B of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0C of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0D of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0E of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0F of ram_2 : label is "4000000000000000000000000000000000000000000000000000000000000000" ;

		attribute INIT_00 of ram_3 : label is "0000000000000343C0F0F030D0CDC0CFF0F00004D4FF00F00000F0DFF4000000" ;
		attribute INIT_01 of ram_3 : label is "208D034D0332D08D034D203384342D08D00F344433444334F310001010001000" ;
		attribute INIT_02 of ram_3 : label is "0F34443034F40030014D4F0401030822003014D4F034D20332033284344DD423" ;
		attribute INIT_03 of ram_3 : label is "35919467843887689804D003D000400300033EC4F0343444E4CE344435583C4F" ;
		attribute INIT_04 of ram_3 : label is "35D0443433421D00F8D03203FF00078003010431D10D110911015910BA431DD4" ;
		attribute INIT_05 of ram_3 : label is "000000000000000000000000000000000000000501030014D4F050000214D4F0" ;
		attribute INIT_06 of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_07 of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_08 of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_09 of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0A of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0B of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0C of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0D of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0E of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0F of ram_3 : label is "1000000000000000000000000000000000000000000000000000000000000000" ;

		attribute INIT_00 of ram_4 : label is "D0A0907070500E4EF00084E00D22000200010202F227F182F2F0400400FF0F00" ;
		attribute INIT_01 of ram_4 : label is "00404D70020000404D60002041E200040000F50FFF50FFF00E40504020E020E0" ;
		attribute INIT_02 of ram_4 : label is "00FB0FFCC00B0C1D004000BA00C1D4104FE0040004D8000200020041E240040E" ;
		attribute INIT_03 of ram_4 : label is "E0C1CF0004EF100380BE00C000DBE0C00D0FF0000C50FC0C01D0FC0FFF3CF300" ;
		attribute INIT_04 of ram_4 : label is "D3004FE0D210000F0400104D0F00000BC2C2D4E10541254122320800784E0004" ;
		attribute INIT_05 of ram_4 : label is "00000000000000000000000000000000000000B500C1D004000B40CD00040004" ;
		attribute INIT_06 of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_07 of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_08 of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_09 of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0A of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0B of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0C of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0D of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0E of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0F of ram_4 : label is "5000000000000000000000000000000000000000000000000000000000000000" ;

		attribute INIT_00 of ram_5 : label is "EEA473C201F000F1F0400F0010900000104F001DF30FD50FEBF000004BD00011" ;
		attribute INIT_01 of ram_5 : label is "12F5FA51100132F4FA811100F030132F40041812E1312F1012DCED1BDAE9485F" ;
		attribute INIT_02 of ram_5 : label is "041A12E00011100721F4015411007F00FF321F401FAB2310011001F030F13F15" ;
		attribute INIT_03 of ram_5 : label is "710707106F67004F01581100107501084701D0001800FF1F1E311812FD08D001" ;
		attribute INIT_04 of ram_5 : label is "AC11F8300002143F4F5000FA0B41004500017F0B3007A003A001F03200F0623F" ;
		attribute INIT_05 of ram_5 : label is "00000000000000000000000000000000000012541100721F40159107321F501F" ;
		attribute INIT_06 of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_07 of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_08 of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_09 of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0A of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0B of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0C of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0D of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0E of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0F of ram_5 : label is "A000000000000000000000000000000000000000000000000000000000000000" ;

		signal data_out : std_logic_vector( 3 downto 0 ) ;
	begin
	    ram_1 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"3131313131310030120203021231020002031313131013131312120003100233",
				INIT_01 => X"0031303112001031303111203100010313202310023100221031313131313131",
				INIT_02 => X"2023100302131303003121331130331031000312130311120112013100311310",
				INIT_03 => X"0313031223031000003311301033313003220002130213131031231001031021",
				INIT_04 => X"0311310110000103131211300000211330333303100330033113310000303113",
				INIT_05 => X"0000000000000000000000000000000000003333113030031213313300031213",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"3000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => data_out,  
				DIB => jdata( JDATASIZE - 1 downto 16 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 
			-- loose top 2 bits
			instruction( 17 downto 16 ) <= data_out( 1 downto 0 ) ;

	    ram_2 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"54545454545460502AAAC40A8F54FA1CCAA54545252A8525454B2A0CA5441C4C",
				INIT_01 => X"6054405C8D76C054405C88D759016C0544AAC5240C524ECB2054545454545454",
				INIT_02 => X"AAC524001B25C0506654B245C80505915206654B2405C88D7C8D78590152C520",
				INIT_03 => X"0545A5C00505400A1645C807C0045C0000AC000B241B45C5C058C5240C154FB2",
				INIT_04 => X"05C8520A91166C05254AFD40DAA6AA8401000505411501150B905466115054C5",
				INIT_05 => X"0000000000000000000000000000000000008045C80706654B245C0066654B24",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"4000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => instruction( 15 downto 12 ),  
				DIB => jdata( 15 downto 12 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 

	    ram_3 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"0000000000000343C0F0F030D0CDC0CFF0F00004D4FF00F00000F0DFF4000000",
				INIT_01 => X"208D034D0332D08D034D203384342D08D00F344433444334F310001010001000",
				INIT_02 => X"0F34443034F40030014D4F0401030822003014D4F034D20332033284344DD423",
				INIT_03 => X"35919467843887689804D003D000400300033EC4F0343444E4CE344435583C4F",
				INIT_04 => X"35D0443433421D00F8D03203FF00078003010431D10D110911015910BA431DD4",
				INIT_05 => X"000000000000000000000000000000000000000501030014D4F050000214D4F0",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"1000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => instruction( 11 downto 8 ),  
				DIB => jdata( 11 downto 8 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 

	    ram_4 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"D0A0907070500E4EF00084E00D22000200010202F227F182F2F0400400FF0F00",
				INIT_01 => X"00404D70020000404D60002041E200040000F50FFF50FFF00E40504020E020E0",
				INIT_02 => X"00FB0FFCC00B0C1D004000BA00C1D4104FE0040004D8000200020041E240040E",
				INIT_03 => X"E0C1CF0004EF100380BE00C000DBE0C00D0FF0000C50FC0C01D0FC0FFF3CF300",
				INIT_04 => X"D3004FE0D210000F0400104D0F00000BC2C2D4E10541254122320800784E0004",
				INIT_05 => X"00000000000000000000000000000000000000B500C1D004000B40CD00040004",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"5000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => instruction( 7 downto 4 ),  
				DIB => jdata( 7 downto 4 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 

	    ram_5 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"EEA473C201F000F1F0400F0010900000104F001DF30FD50FEBF000004BD00011",
				INIT_01 => X"12F5FA51100132F4FA811100F030132F40041812E1312F1012DCED1BDAE9485F",
				INIT_02 => X"041A12E00011100721F4015411007F00FF321F401FAB2310011001F030F13F15",
				INIT_03 => X"710707106F67004F01581100107501084701D0001800FF1F1E311812FD08D001",
				INIT_04 => X"AC11F8300002143F4F5000FA0B41004500017F0B3007A003A001F03200F0623F",
				INIT_05 => X"00000000000000000000000000000000000012541100721F40159107321F501F",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"A000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => instruction( 3 downto 0 ),  
				DIB => jdata( 3 downto 0 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 
	end generate ;

	jdata <= ( others => '0' ) ;
	jaddr <= ( others => '0' ) ;
	juser1 <= '0' ;
	jwrite <= '0' ;
end architecture mix ;

